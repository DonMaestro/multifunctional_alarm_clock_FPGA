

module testing_block(display_bus A);




endmodule
